package some_package;
    parameter foo = 0;
endpackage : some_package